`default_nettype none

module snitch_logo ();
endmodule
