VERSION 5.8 ;

MACRO snitch_names_small_logo
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN snitch_small_logo 0 0 ;
  SIZE 150 BY 150 ;

  OBS
    LAYER TopMetal1 ;
      RECT 0 0 150 150 ;
  END
END snitch_small_logo
