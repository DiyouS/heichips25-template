`default_nettype none

module snitch_names_small_logo ();
endmodule
